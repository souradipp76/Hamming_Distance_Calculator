* SPICE NETLIST
***************************************

.SUBCKT nwell_contact
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT fuladdlay Cin IN1 IN2 S VDD GND Cout
** N=18 EP=7 IP=5 FDC=30
M0 S 3 6 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-24200 $Y=-44250 $D=1
M1 3 IN2 7 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-23950 $Y=-12300 $D=1
M2 3 6 S GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-850 $Y=-44350 $D=1
M3 IN2 7 3 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-600 $Y=-12200 $D=1
M4 GND Cin 6 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=22150 $Y=-44250 $D=1
M5 GND IN1 7 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=22400 $Y=-12300 $D=1
M6 10 Cin 8 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=44300 $Y=-44200 $D=1
M7 11 IN1 9 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=44550 $Y=-12350 $D=1
M8 GND 3 8 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=66350 $Y=-44100 $D=1
M9 GND IN2 9 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=66600 $Y=-12450 $D=1
M10 5 10 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=88650 $Y=-44050 $D=1
M11 15 11 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=88900 $Y=-12500 $D=1
M12 GND 15 12 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=111100 $Y=-12550 $D=1
M13 12 5 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=134500 $Y=-12600 $D=1
M14 Cout 12 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=157400 $Y=-12600 $D=1
M15 S 3 Cin VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-24200 $Y=-71600 $D=0
M16 3 IN2 IN1 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-23950 $Y=5050 $D=0
M17 3 Cin S VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-850 $Y=-71700 $D=0
M18 IN2 IN1 3 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-600 $Y=5150 $D=0
M19 VDD Cin 6 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=22150 $Y=-71600 $D=0
M20 VDD IN1 7 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=22400 $Y=5050 $D=0
M21 10 Cin VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=44300 $Y=-71550 $D=0
M22 11 IN1 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=44550 $Y=5000 $D=0
M23 VDD 3 10 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=66350 $Y=-71450 $D=0
M24 VDD IN2 11 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=66600 $Y=4900 $D=0
M25 5 10 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=88650 $Y=-71400 $D=0
M26 15 11 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=88900 $Y=4850 $D=0
M27 16 15 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=111100 $Y=4800 $D=0
M28 12 5 16 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=134500 $Y=4750 $D=0
M29 Cout 12 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=157400 $Y=4750 $D=0
.ENDS
***************************************

* ELDO netlist generated with ICnet by 'vlsi' on Fri Oct 20 2017 at 02:29:08

.CONNECT GND 0

*
* Component pathname : /home/vlsi/dff/inverter.cir
*
.subckt INVERTER_CIR_ESC1  OUT GND IN VDD

        MN1 OUT IN GND VSS n L=1.8e-07 W=1.9e-07
        MP1 OUT IN VDD VDD p L=1.8e-07 W=1.31e-06
.ends INVERTER_CIR_ESC1

*
* Component pathname : /home/vlsi/dff/Dflipflopnoinvnew.cir
*
.subckt DFLIPFLOPNOINVNEW_CIR_ESC2  OUT CLK D GND NCLK VDD

        MN2 N$7 CLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP2 N$7 NCLK N$56 VDD p L=1.8e-07 W=1.31e-06
        MN1 N$4 NCLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP1 N$4 CLK N$56 VDD p L=1.8e-07 W=1.31e-06
        X_INVERTER_CIR3_ESC3 OUT GND N$56 VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR2_ESC4 N$7 GND D VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR1_ESC5 N$4 GND OUT VDD INVERTER_CIR_ESC1
.ends DFLIPFLOPNOINVNEW_CIR_ESC2

*
* Component pathname : /home/vlsi/dff/masterslaveDflipflopnew.cir
*
.subckt MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6  OUT CLEAR CLK D GND NCLK PRESET
+ VDD

        X_DFLIPFLOPNOINVNEW_CIR1_ESC7 N$34 NCLK D GND CLK VDD DFLIPFLOPNOINVNEW_CIR_ESC2
        X_DFLIPFLOPNOINVNEW_CIR2_ESC8 OUT CLK N$34 GND NCLK VDD DFLIPFLOPNOINVNEW_CIR_ESC2
.ends MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6

*
* Component pathname : /home/vlsi/g4/or
*
.subckt OR  OUT GND IN1 IN2 VDD

        MN3 OUT N$7 GND VSS n L=1.8e-07 W=3.6e-07
        MP3 OUT N$7 VDD VDD p L=1.8e-07 W=1.26e-06
        MN2 N$7 IN2 GND VSS n L=1.8e-07 W=3.6e-07
        MN1 N$7 IN1 GND VSS n L=1.8e-07 W=3.6e-07
        MP2 N$5 IN1 VDD VDD p L=1.8e-07 W=2.52e-06
        MP1 N$7 IN2 N$5 VDD p L=1.8e-07 W=2.52e-06
.ends OR

*
* Component pathname : /home/vlsi/g4/xor
*
.subckt XOR  OUT GND IN1 IN2 VDD

        MN7 OUT N$22 GND VSS n L=1.8e-07 W=3.6e-07
        MP7 OUT N$22 VDD VDD p L=1.8e-07 W=1.26e-06
        MP6 N$47 IN2 VDD VDD p L=1.8e-07 W=1.26e-06
        MN6 N$47 IN2 GND VSS n L=1.8e-07 W=3.6e-07
        MP5 N$59 IN1 VDD VDD p L=1.8e-07 W=1.26e-06
        MN5 N$59 IN1 GND VSS n L=1.8e-07 W=3.6e-07
        MN1 N$22 N$59 N$24 VSS n L=1.8e-07 W=7.2e-07
        MN4 N$2 N$47 GND VSS n L=1.8e-07 W=7.2e-07
        MN3 N$24 IN2 GND VSS n L=1.8e-07 W=7.2e-07
        MN2 N$22 IN1 N$2 VSS n L=1.8e-07 W=7.2e-07
        MP4 N$22 N$47 N$7 VDD p L=1.8e-07 W=2.52e-06
        MP3 N$7 N$59 VDD VDD p L=1.8e-07 W=2.52e-06
        MP2 N$22 IN2 N$31 VDD p L=1.8e-07 W=2.52e-06
        MP1 N$31 IN1 VDD VDD p L=1.8e-07 W=2.52e-06
.ends XOR

*
* Component pathname : /home/vlsi/g4/and
*
.subckt AND  OUT GND IN1 IN2 VDD

        MP3 OUT N$5 VDD VDD p L=1.8e-07 W=1.26e-06
        MN3 OUT N$5 GND VSS n L=1.8e-07 W=3.6e-07
        MP2 N$5 IN2 VDD VDD p L=1.8e-07 W=1.26e-06
        MP1 N$5 IN1 VDD VDD p L=1.8e-07 W=1.26e-06
        MN2 N$2 IN2 GND VSS n L=1.8e-07 W=7.2e-07
        MN1 N$5 IN1 N$2 VSS n L=1.8e-07 W=7.2e-07
.ends AND

*
* Component pathname : /home/vlsi/g4/halfadd
*
.subckt HALFADD  C S GND IN1 IN2 VDD

        X_EXC1 S GND IN1 IN2 VDD XOR
        X_AND1 C GND IN2 IN1 VDD AND
.ends HALFADD

*
* Component pathname : /home/vlsi/g4/fulladd
*
.subckt FULLADD  C S CIN GND IN1 IN2 VDD

        X_OR1 C GND N$16 N$13 VDD OR
        X_HALFADD2 N$16 S GND N$11 CIN VDD HALFADD
        X_HALFADD1 N$13 N$11 GND IN2 IN1 VDD HALFADD
.ends FULLADD

*
* Component pathname : /home/vlsi/dff/mux.cir
*
.subckt MUX_CIR_ESC9  OUT GND IN1 IN2 S VDD

        MN3 N$3 S GND VSS n L=1.8e-07 W=3.6e-07
        MP3 N$3 S VDD VDD p L=1.8e-07 W=1.26e-06
        MN2 IN2 N$3 OUT VSS n L=1.8e-07 W=3.6e-07
        MP2 IN2 S OUT VDD p L=1.8e-07 W=1.26e-06
        MN1 IN1 S OUT VSS n L=1.8e-07 W=3.6e-07
        MP1 IN1 N$3 OUT VDD p L=1.8e-07 W=1.26e-06
.ends MUX_CIR_ESC9

*
* Component pathname : /home/vlsi/dff/sipopisonew.cir
*
.subckt SIPOPISONEW_CIR_ESC10  P1 P2 P3 CLK GND L1 L2 L3 NCLK SEL SIN VDD

        X_MUX_CIR3_ESC11 N$14 GND L3 P2 SEL VDD MUX_CIR_ESC9
        X_MUX_CIR2_ESC12 N$10 GND L2 P1 SEL VDD MUX_CIR_ESC9
        X_MUX_CIR1_ESC13 N$3 GND L1 SIN SEL VDD MUX_CIR_ESC9
        X_Q3 P3 N$13 CLK N$14 GND NCLK N$16 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_Q2 P2 N$9 CLK N$10 GND NCLK N$12 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_Q1 P1 N$1 CLK N$3 GND NCLK N$7 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
.ends SIPOPISONEW_CIR_ESC10

*
* MAIN CELL: Component pathname : /home/vlsi/g4/multi
*
        X_MASTERSLAVEDFLIPFLOPNEW_CIR10_ESC14 N$91 N$149 CLK N$89 GND NCLK
+ N$150 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_MASTERSLAVEDFLIPFLOPNEW_CIR6_ESC15 N$78 N$147 CLK N$76 GND NCLK
+ N$148 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_FULLADD2 N$89 N$92 N$91 GND N$83 N$87 VDD FULLADD
        X_FULLADD1 N$76 N$83 N$78 GND N$80 N$74 VDD FULLADD
        X_AND3 N$87 GND IN N$64 VDD AND
        X_AND2 N$80 GND IN N$61 VDD AND
        X_AND1 N$74 GND IN N$58 VDD AND
        X_MASTERSLAVEDFLIPFLOPNEW_CIR8_ESC16 O4 N$21 CLK O3 GND NCLK N$52
+ VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_MASTERSLAVEDFLIPFLOPNEW_CIR7_ESC17 O3 N$16 CLK O2 GND NCLK N$49
+ VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_MASTERSLAVEDFLIPFLOPNEW_CIR9_ESC18 O5 N$26 CLK O4 GND NCLK N$55
+ VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_MASTERSLAVEDFLIPFLOPNEW_CIR5_ESC19 O2 N$11 CLK O1 GND NCLK N$46
+ VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_MASTERSLAVEDFLIPFLOPNEW_CIR4_ESC20 O1 N$6 CLK O0 GND NCLK N$43
+ VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_MASTERSLAVEDFLIPFLOPNEW_CIR3_ESC21 O0 N$1 CLK N$92 GND NCLK N$40
+ VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_MASTERSLAVEDFLIPFLOPNEW_CIR2_ESC22 N$64 N$145 CLK N$61 GND NCLK
+ N$146 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_MASTERSLAVEDFLIPFLOPNEW_CIR1_ESC23 N$61 N$143 CLK N$58 GND NCLK
+ N$144 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_SIPOPISONEW_CIR1_ESC24 N$139 N$140 N$58 CLK GND IN IN IN NCLK
+ SEL IN VDD SIPOPISONEW_CIR_ESC10
*
.end

* SPICE NETLIST
***************************************

.SUBCKT nwell_contact
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT dhallsipolay in clk ~clk out3 out1 out2 gnd vdd
** N=29 EP=8 IP=2 FDC=60
M0 13 in gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=157550 $Y=-5850 $D=1
M1 14 out1 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=157850 $Y=-42900 $D=1
M2 15 out2 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=158050 $Y=-152250 $D=1
M3 7 ~clk 13 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=179650 $Y=-5850 $D=1
M4 8 ~clk 14 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=179950 $Y=-42900 $D=1
M5 9 ~clk 15 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=180150 $Y=-152250 $D=1
M6 7 clk 16 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=204200 $Y=-5950 $D=1
M7 8 clk 17 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=204500 $Y=-42800 $D=1
M8 9 clk 18 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=204700 $Y=-152350 $D=1
M9 19 7 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=226250 $Y=-6000 $D=1
M10 20 8 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=226550 $Y=-42750 $D=1
M11 21 9 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=226750 $Y=-152400 $D=1
M12 16 19 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=248500 $Y=-6000 $D=1
M13 17 20 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=248800 $Y=-42750 $D=1
M14 18 21 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=249000 $Y=-152400 $D=1
M15 22 19 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=270750 $Y=-6000 $D=1
M16 23 20 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=271050 $Y=-42750 $D=1
M17 24 21 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=271250 $Y=-152400 $D=1
M18 10 clk 22 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=292850 $Y=-6000 $D=1
M19 11 clk 23 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=293150 $Y=-42750 $D=1
M20 12 clk 24 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=293350 $Y=-152400 $D=1
M21 10 ~clk 25 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=317400 $Y=-6100 $D=1
M22 11 ~clk 26 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=317700 $Y=-42650 $D=1
M23 12 ~clk 27 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=317900 $Y=-152500 $D=1
M24 out1 10 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=339450 $Y=-6150 $D=1
M25 out2 11 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=339750 $Y=-42600 $D=1
M26 out3 12 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=339950 $Y=-152550 $D=1
M27 25 out1 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=361700 $Y=-6150 $D=1
M28 26 out2 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=362000 $Y=-42600 $D=1
M29 27 out3 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=362200 $Y=-152550 $D=1
M30 13 in vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=157550 $Y=15550 $D=0
M31 14 out1 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=157850 $Y=-74300 $D=0
M32 15 out2 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=158050 $Y=-130850 $D=0
M33 7 ~clk 16 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=179650 $Y=15550 $D=0
M34 8 ~clk 17 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=179950 $Y=-74300 $D=0
M35 9 ~clk 18 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=180150 $Y=-130850 $D=0
M36 7 clk 13 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=204200 $Y=15450 $D=0
M37 8 clk 14 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=204500 $Y=-74200 $D=0
M38 9 clk 15 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=204700 $Y=-130950 $D=0
M39 19 7 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=226250 $Y=15400 $D=0
M40 20 8 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=226550 $Y=-74150 $D=0
M41 21 9 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=226750 $Y=-131000 $D=0
M42 16 19 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=248500 $Y=15400 $D=0
M43 17 20 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=248800 $Y=-74150 $D=0
M44 18 21 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=249000 $Y=-131000 $D=0
M45 22 19 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=270750 $Y=15400 $D=0
M46 23 20 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=271050 $Y=-74150 $D=0
M47 24 21 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=271250 $Y=-131000 $D=0
M48 10 clk 25 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=292850 $Y=15400 $D=0
M49 11 clk 26 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=293150 $Y=-74150 $D=0
M50 12 clk 27 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=293350 $Y=-131000 $D=0
M51 10 ~clk 22 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=317400 $Y=15300 $D=0
M52 11 ~clk 23 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=317700 $Y=-74050 $D=0
M53 12 ~clk 24 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=317900 $Y=-131100 $D=0
M54 out1 10 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=339450 $Y=15250 $D=0
M55 out2 11 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=339750 $Y=-74000 $D=0
M56 out3 12 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=339950 $Y=-131150 $D=0
M57 25 out1 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=361700 $Y=15250 $D=0
M58 26 out2 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=362000 $Y=-74000 $D=0
M59 27 out3 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=362200 $Y=-131150 $D=0
.ENDS
***************************************

* ELDO netlist generated with ICnet by 'vlsi' on Sun Oct 29 2017 at 23:10:28

.CONNECT GND 0

*
* MAIN CELL: Component pathname : /home/vlsi/g4/exc
*
        MP4 OUT IN1 IN2 VDD p L=1.8e-07 W=1.26e-06
        MN4 OUT N$32 IN2 VSS n L=1.8e-07 W=3.6e-07
        MN2 N$32 IN1 GND VSS n L=1.8e-07 W=3.6e-07
        MP2 N$32 IN1 VDD VDD p L=1.8e-07 W=1.26e-06
        MN1 OUT IN2 N$32 VSS n L=1.8e-07 W=3.6e-07
        MP1 OUT IN2 IN1 VDD p L=1.8e-07 W=1.26e-06
*
.end

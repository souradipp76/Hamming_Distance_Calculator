* ELDO netlist generated with ICnet by 'vlsi' on Thu Oct 19 2017 at 00:44:36

.CONNECT GND 0

*
* Component pathname : /home/vlsi/dff/mux.cir
*
.subckt MUX_CIR_ESC1  OUT GND IN1 IN2 S VDD

        MN3 N$3 S GND VSS n L=1.8e-07 W=3.6e-07
        MP3 N$3 S VDD VDD p L=1.8e-07 W=1.26e-06
        MN2 IN2 N$3 OUT VSS n L=1.8e-07 W=3.6e-07
        MP2 IN2 S OUT VDD p L=1.8e-07 W=1.26e-06
        MN1 IN1 S OUT VSS n L=1.8e-07 W=3.6e-07
        MP1 IN1 N$3 OUT VDD p L=1.8e-07 W=1.26e-06
.ends MUX_CIR_ESC1

*
* Component pathname : /home/vlsi/dff/inverter.cir
*
.subckt INVERTER_CIR_ESC2  OUT GND IN VDD

        MN1 OUT IN GND VSS n L=1.8e-07 W=1.9e-07
        MP1 OUT IN VDD VDD p L=1.8e-07 W=1.31e-06
.ends INVERTER_CIR_ESC2

*
* Component pathname : /home/vlsi/dff/Dflipflopnoinvnew.cir
*
.subckt DFLIPFLOPNOINVNEW_CIR_ESC3  OUT CLK D GND NCLK VDD

        MN2 N$7 CLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP2 N$7 NCLK N$56 VDD p L=1.8e-07 W=1.31e-06
        MN1 N$4 NCLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP1 N$4 CLK N$56 VDD p L=1.8e-07 W=1.31e-06
        X_INVERTER_CIR3_ESC4 OUT GND N$56 VDD INVERTER_CIR_ESC2
        X_INVERTER_CIR2_ESC5 N$7 GND D VDD INVERTER_CIR_ESC2
        X_INVERTER_CIR1_ESC6 N$4 GND OUT VDD INVERTER_CIR_ESC2
.ends DFLIPFLOPNOINVNEW_CIR_ESC3

*
* Component pathname : /home/vlsi/dff/masterslaveDflipflopnew.cir
*
.subckt MASTERSLAVEDFLIPFLOPNEW_CIR_ESC7  OUT CLEAR CLK D GND NCLK PRESET
+ VDD

        X_DFLIPFLOPNOINVNEW_CIR1_ESC8 N$34 NCLK D GND CLK VDD DFLIPFLOPNOINVNEW_CIR_ESC3
        X_DFLIPFLOPNOINVNEW_CIR2_ESC9 OUT CLK N$34 GND NCLK VDD DFLIPFLOPNOINVNEW_CIR_ESC3
.ends MASTERSLAVEDFLIPFLOPNEW_CIR_ESC7

*
* MAIN CELL: Component pathname : /home/vlsi/g4/serdes
*
        X_MUX_CIR3_ESC10 N$14 GND L3 P2 SEL VDD MUX_CIR_ESC1
        X_MUX_CIR2_ESC11 N$10 GND L2 P1 SEL VDD MUX_CIR_ESC1
        X_MUX_CIR1_ESC12 N$3 GND L1 SIN SEL VDD MUX_CIR_ESC1
        X_Q3 P3 N$13 CLK N$14 GND NCLK N$16 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC7
        X_Q2 P2 N$9 CLK N$10 GND NCLK N$12 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC7
        X_Q1 P1 N$1 CLK N$3 GND NCLK N$7 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC7
*
.end

* Component: /home/vlsi/g4/halfadd Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/halfadd/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0 100n 0

* --- Forces
VFORCE__GND GND GND DC 0
VFORCE__VDD VDD GND DC 1.8
VFORCE__IN1 IN1 GND PULSE (0 1 0 1n 1n 20n 50n)
VFORCE__IN2 IN2 GND PULSE (0 1 0 1n 1n 10n 25n)

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT TRAN V(S) V(IN1) V(C) V(IN2)

* --- Params
.TEMP 27.0

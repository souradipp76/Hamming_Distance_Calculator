* Component: /home/vlsi/dff/mux.cir Viewpoint: tsmc018a

.INCLUDE /home/vlsi/dff/mux.cir/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0 100n 0 UIC

* --- Forces
VFORCE__GND GND GND DC 0
VFORCE__VDD VDD GND DC 1.8
VFORCE__IN1 IN1 GND PULSE (0 1.8 0u 1n 1n 10n 25n)
VFORCE__IN2 IN2 GND PULSE (0 1.8 0u 1n 1n 20n 50n)
VFORCE__S S GND PULSE (0 1.8 0u 1n 1n 30n 60n)

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PROBE TRAN V(OUT)

* --- Params
.TEMP 27.0

* SPICE NETLIST
***************************************

.SUBCKT answer_lay D CLK_INV CLK Out Vdd Gnd
** N=13 EP=6 IP=0 FDC=20
M0 7 D Gnd Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-6900 $Y=-45400 $D=1
M1 2 CLK_INV 7 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=47250 $Y=-46300 $D=1
M2 8 CLK 2 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=112500 $Y=-47600 $D=1
M3 Gnd 9 8 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=166650 $Y=-48500 $D=1
M4 Gnd 2 9 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=228550 $Y=-49150 $D=1
M5 10 9 Gnd Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=337750 $Y=-51000 $D=1
M6 5 CLK 10 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=391900 $Y=-51900 $D=1
M7 11 CLK_INV 5 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=457150 $Y=-53200 $D=1
M8 Gnd Out 11 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=511300 $Y=-54100 $D=1
M9 Gnd 5 Out Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=573200 $Y=-54750 $D=1
M10 7 D Vdd Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-6900 $Y=5500 $D=0
M11 2 CLK 7 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=47250 $Y=4600 $D=0
M12 8 CLK_INV 2 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=112500 $Y=3300 $D=0
M13 Vdd 9 8 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=166650 $Y=2400 $D=0
M14 Vdd 2 9 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=228550 $Y=1750 $D=0
M15 10 9 Vdd Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=337750 $Y=-100 $D=0
M16 5 CLK_INV 10 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=391900 $Y=-1000 $D=0
M17 11 CLK 5 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=457150 $Y=-2300 $D=0
M18 Vdd Out 11 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=511300 $Y=-3200 $D=0
M19 Vdd 5 Out Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=573200 $Y=-3850 $D=0
.ENDS
***************************************

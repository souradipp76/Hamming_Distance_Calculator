* Component: /home/vlsi/g4/sipo.cir Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/sipo.cir/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - DCOP
.OPTION PROBEOP2
.OP

* - Analysis Setup - Trans
.TRAN 0 300n 0 UIC

* --- Forces
VFORCE__GND GND GND DC 0
VFORCE__VDD VDD GND DC 1.8
VFORCE__CLK CLK GND PULSE (0 1.8 5n 1n 1n 20n 50n)
VFORCE__NCLK NCLK GND PULSE (1.8 0 5n 1n 1n 20n 50n)
VFORCE__SIN SIN GND PATTERN 5 0 0 1n 1n 50n 11011 R=0.0

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT DC V(P3) V(P2) V(P1)
.PLOT TRAN V(P3) V(P2) V(P1)

* --- Params
.TEMP 27.0

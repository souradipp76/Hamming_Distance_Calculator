* Component: /home/vlsi/g4/exc Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/exc/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0 150n 0

* --- Forces
VFORCE__VDD VDD GND DC 1.8
VFORCE__GND GND GND DC 0
VFORCE__IN1 IN1 GND PATTERN 1.8 0 0 1n 1n 50n 000 R=0.0
VFORCE__IN2 IN2 GND PATTERN 1.8 0 0 1n 1n 50n 111 R=0.0

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT TRAN V(IN1) V(IN2) V(OUT)

* --- Params
.TEMP 27.0

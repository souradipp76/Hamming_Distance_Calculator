* ELDO netlist generated with ICnet by 'vlsi' on Tue Oct  3 2017 at 10:13:16

.CONNECT GND 0

*
* Component pathname : /home/vlsi/dff/inverter.cir
*
.subckt INVERTER_CIR_ESC1  OUT GND IN VDD

        MN1 OUT IN GND VSS n L=1.8e-07 W=1.9e-07
        MP1 OUT IN VDD VDD p L=1.8e-07 W=1.31e-06
.ends INVERTER_CIR_ESC1

*
* MAIN CELL: Component pathname : /home/vlsi/dff/Dflipflopnoinvnew.cir
*
        MN2 N$7 CLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP2 N$7 NCLK N$56 VDD p L=1.8e-07 W=1.31e-06
        MN1 N$4 NCLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP1 N$4 CLK N$56 VDD p L=1.8e-07 W=1.31e-06
        X_INVERTER_CIR3_ESC2 OUT GND N$56 VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR2_ESC3 N$7 GND D VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR1_ESC4 N$4 GND OUT VDD INVERTER_CIR_ESC1
*
.end

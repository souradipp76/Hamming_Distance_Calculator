* Component: /home/vlsi/g4/dhall_flip Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/dhall_flip/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - DCOP
.OPTION PROBEOP2
.OP

* - Analysis Setup - Trans
.TRAN 0.0 100n 0

* --- Forces
VFORCE___VDD VDD GND DC 1.8
VFORCE___GND GND GND DC 0
VFORCE__D D GND DC 1.8
VFORCE__~clk N_CLK_ESC1 GND PULSE (1.8 0 5n 1n 1n 20n 50n)
VFORCE__clk CLK GND PULSE (0 1.8 5n 1n 1n 20n 50n)

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT DC V(OUT)
.PLOT TRAN V(OUT)

* --- Params
.TEMP 27.0

* ELDO netlist generated with ICnet by 'vlsi' on Thu Oct 19 2017 at 00:57:11

.CONNECT GND 0

*
* Component pathname : /home/vlsi/g4/xor
*
.subckt XOR  OUT GND IN1 IN2 VDD

        MN7 OUT N$22 GND VSS n L=1.8e-07 W=3.6e-07
        MP7 OUT N$22 VDD VDD p L=1.8e-07 W=1.26e-06
        MP6 N$47 IN2 VDD VDD p L=1.8e-07 W=1.26e-06
        MN6 N$47 IN2 GND VSS n L=1.8e-07 W=3.6e-07
        MP5 N$59 IN1 VDD VDD p L=1.8e-07 W=1.26e-06
        MN5 N$59 IN1 GND VSS n L=1.8e-07 W=3.6e-07
        MN1 N$22 N$59 N$24 VSS n L=1.8e-07 W=7.2e-07
        MN4 N$2 N$47 GND VSS n L=1.8e-07 W=7.2e-07
        MN3 N$24 IN2 GND VSS n L=1.8e-07 W=7.2e-07
        MN2 N$22 IN1 N$2 VSS n L=1.8e-07 W=7.2e-07
        MP4 N$22 N$47 N$7 VDD p L=1.8e-07 W=2.52e-06
        MP3 N$7 N$59 VDD VDD p L=1.8e-07 W=2.52e-06
        MP2 N$22 IN2 N$31 VDD p L=1.8e-07 W=2.52e-06
        MP1 N$31 IN1 VDD VDD p L=1.8e-07 W=2.52e-06
.ends XOR

*
* Component pathname : /home/vlsi/g4/and
*
.subckt AND  OUT GND IN1 IN2 VDD

        MP3 OUT N$5 VDD VDD p L=1.8e-07 W=1.26e-06
        MN3 OUT N$5 GND VSS n L=1.8e-07 W=3.6e-07
        MP2 N$5 IN2 VDD VDD p L=1.8e-07 W=1.26e-06
        MP1 N$5 IN1 VDD VDD p L=1.8e-07 W=1.26e-06
        MN2 N$2 IN2 GND VSS n L=1.8e-07 W=7.2e-07
        MN1 N$5 IN1 N$2 VSS n L=1.8e-07 W=7.2e-07
.ends AND

*
* MAIN CELL: Component pathname : /home/vlsi/g4/halfadd
*
        X_EXC1 S GND IN1 IN2 VDD XOR
        X_AND1 C GND IN2 IN1 VDD AND
*
.end

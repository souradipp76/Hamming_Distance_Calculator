* Component: /home/vlsi/g4/dhall_sipo Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/dhall_sipo/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0 150n 0

* --- Forces
VFORCE__clk CLK GND PULSE (0 1.8 15n 1n 1n 20n 50n)
VFORCE__GND_1 GND GND DC 0
VFORCE__VDD VDD GND DC 1.8
VFORCE__IN1 IN1 GND PATTERN 1.8 0 0 1n 1n 50n 101 R=0.0
VFORCE__IN2 IN2 GND PATTERN 1.8 0 0 1n 1n 50n 001 R=0.0

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT TRAN V(S1) V(S0)

* --- Params
.TEMP 27.0

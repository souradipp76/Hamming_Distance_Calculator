* File: dhallsipolay_pex.sp
* Created: Sat Oct 28 12:27:26 2017
* Program "Calibre xRC"
* Version "v2013.4_37.29"
* 
.include "dhallsipolay_pex.sp.pex"
.subckt DHALLSIPOLAY  IN CLK :CLK OUT3 OUT1 OUT2 GND VDD
* 
* VDD	VDD
* GND	GND
* OUT2	OUT2
* OUT1	OUT1
* OUT3	OUT3
* ~CLK	~CLK
* CLK	CLK
* IN	IN
M0 N_13_M0_d N_IN_M0_g N_GND_M0_s N_GND_M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M1 N_14_M1_d N_OUT1_M1_g N_GND_M1_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M2 N_15_M2_d N_OUT2_M2_g N_GND_M2_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M3 N_7_M3_d N_:CLK_M3_g N_13_M3_s N_GND_M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M4 N_8_M4_d N_:CLK_M4_g N_14_M4_s N_GND_M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M5 N_9_M5_d N_:CLK_M5_g N_15_M5_s N_GND_M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M6 N_7_M6_d N_CLK_M6_g N_16_M6_s N_GND_M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M7 N_8_M7_d N_CLK_M7_g N_17_M7_s N_GND_M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M8 N_9_M8_d N_CLK_M8_g N_18_M8_s N_GND_M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M9 N_19_M9_d N_7_M9_g N_GND_M9_s N_GND_M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M10 N_20_M10_d N_8_M10_g N_GND_M10_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M11 N_21_M11_d N_9_M11_g N_GND_M11_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M12 N_16_M12_d N_19_M12_g N_GND_M12_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M13 N_17_M13_d N_20_M13_g N_GND_M13_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M14 N_18_M14_d N_21_M14_g N_GND_M14_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M15 N_22_M15_d N_19_M15_g N_GND_M15_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M16 N_23_M16_d N_20_M16_g N_GND_M16_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M17 N_24_M17_d N_21_M17_g N_GND_M17_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M18 N_10_M18_d N_CLK_M18_g N_22_M18_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M19 N_11_M19_d N_CLK_M19_g N_23_M19_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M20 N_12_M20_d N_CLK_M20_g N_24_M20_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M21 N_10_M21_d N_:CLK_M21_g N_25_M21_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M22 N_11_M22_d N_:CLK_M22_g N_26_M22_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M23 N_12_M23_d N_:CLK_M23_g N_27_M23_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M24 N_OUT1_M24_d N_10_M24_g N_GND_M24_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M25 N_OUT2_M25_d N_11_M25_g N_GND_M25_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M26 N_OUT3_M26_d N_12_M26_g N_GND_M26_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M27 N_25_M27_d N_OUT1_M27_g N_GND_M27_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M28 N_26_M28_d N_OUT2_M28_g N_GND_M28_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M29 N_27_M29_d N_OUT3_M29_g N_GND_M29_s N_GND_M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M30 N_13_M30_d N_IN_M30_g N_VDD_M30_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M31 N_14_M31_d N_OUT1_M31_g N_VDD_M31_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M32 N_15_M32_d N_OUT2_M32_g N_VDD_M32_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M33 N_7_M33_d N_:CLK_M33_g N_16_M33_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M34 N_8_M34_d N_:CLK_M34_g N_17_M34_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M35 N_9_M35_d N_:CLK_M35_g N_18_M35_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M36 N_7_M36_d N_CLK_M36_g N_13_M36_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M37 N_8_M37_d N_CLK_M37_g N_14_M37_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M38 N_9_M38_d N_CLK_M38_g N_15_M38_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M39 N_19_M39_d N_7_M39_g N_VDD_M39_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M40 N_20_M40_d N_8_M40_g N_VDD_M40_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M41 N_21_M41_d N_9_M41_g N_VDD_M41_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M42 N_16_M42_d N_19_M42_g N_VDD_M42_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M43 N_17_M43_d N_20_M43_g N_VDD_M43_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M44 N_18_M44_d N_21_M44_g N_VDD_M44_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M45 N_22_M45_d N_19_M45_g N_VDD_M45_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M46 N_23_M46_d N_20_M46_g N_VDD_M46_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M47 N_24_M47_d N_21_M47_g N_VDD_M47_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M48 N_10_M48_d N_CLK_M48_g N_25_M48_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M49 N_11_M49_d N_CLK_M49_g N_26_M49_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M50 N_12_M50_d N_CLK_M50_g N_27_M50_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M51 N_10_M51_d N_:CLK_M51_g N_22_M51_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M52 N_11_M52_d N_:CLK_M52_g N_23_M52_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M53 N_12_M53_d N_:CLK_M53_g N_24_M53_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M54 N_OUT1_M54_d N_10_M54_g N_VDD_M54_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M55 N_OUT2_M55_d N_11_M55_g N_VDD_M55_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M56 N_OUT3_M56_d N_12_M56_g N_VDD_M56_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M57 N_25_M57_d N_OUT1_M57_g N_VDD_M57_s N_VDD_M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M58 N_26_M58_d N_OUT2_M58_g N_VDD_M58_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M59 N_27_M59_d N_OUT3_M59_g N_VDD_M59_s N_VDD_M31_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
*
.include "dhallsipolay_pex.sp.DHALLSIPOLAY.pxi"
*
.ends
*
*

* ELDO netlist generated with ICnet by 'vlsi' on Tue Oct 10 2017 at 11:27:22

.CONNECT GND 0


*
* Component pathname : /home/vlsi/mux [SPICE]
*
*       .include /home/vlsi/mux/asim_lib/mux

*
* Component pathname : /home/vlsi/dff/inverter.cir
*
.subckt INVERTER_CIR_ESC1  OUT GND IN VDD

        MN1 OUT IN GND VSS n L=1.8e-07 W=1.9e-07
        MP1 OUT IN VDD VDD p L=1.8e-07 W=1.31e-06
.ends INVERTER_CIR_ESC1

*
* Component pathname : /home/vlsi/dff/Dflipflopnoinvnew.cir
*
.subckt DFLIPFLOPNOINVNEW_CIR_ESC2  OUT CLK D GND NCLK VDD

        MN2 N$7 CLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP2 N$7 NCLK N$56 VDD p L=1.8e-07 W=1.31e-06
        MN1 N$4 NCLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP1 N$4 CLK N$56 VDD p L=1.8e-07 W=1.31e-06
        X_INVERTER_CIR3_ESC3 OUT GND N$56 VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR2_ESC4 N$7 GND D VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR1_ESC5 N$4 GND OUT VDD INVERTER_CIR_ESC1
.ends DFLIPFLOPNOINVNEW_CIR_ESC2

*
* Component pathname : /home/vlsi/dff/masterslaveDflipflopnew.cir
*
.subckt MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6  OUT CLK D GND NCLK VDD

        X_DFLIPFLOPNOINVNEW_CIR1_ESC7 N$34 NCLK D GND CLK VDD DFLIPFLOPNOINVNEW_CIR_ESC2
        X_DFLIPFLOPNOINVNEW_CIR2_ESC8 OUT CLK N$34 GND NCLK VDD DFLIPFLOPNOINVNEW_CIR_ESC2
.ends MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6

*
* MAIN CELL: Component pathname : /home/vlsi/dff/sipopiso.cir
*
        X_MUX3 N$83 GND D PO3 S VDD mux
        X_MUX2 N$82 GND C PO2 S VDD mux
        X_MUX1 N$81 GND B PO1 S VDD mux
        X_MUX5 N$80 GND A SIN S VDD mux
        X_I$5 N$27 GND CLK VDD INVERTER_CIR_ESC1
        X_I$4 SO CLK N$83 GND N$27 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_I$3 PO3 CLK N$82 GND N$27 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_I$2 PO2 CLK N$81 GND N$27 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_I$1 PO1 CLK N$80 GND N$27 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
*
.end

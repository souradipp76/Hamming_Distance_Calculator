* Component: /home/vlsi/g4/or Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/or/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0 100n 0

* --- Forces
VFORCE__GND VDD GND DC 1.8
VFORCE__GND_1 GND GND DC 0
VFORCE__IN2 IN2 GND PULSE (0 1.8 0 1n 1n 10n 25n)
VFORCE__IN1_1 IN1 GND PULSE (0 1.8 0 1n 1n 20n 50n)

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT TRAN V(OUT) V(IN2) V(IN1)

* --- Params
.TEMP 27

* Component: /home/vlsi/g4/faddfinal Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/faddfinal/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0 100n 0

* --- Forces
VFORCE__Cin IN1 GND DC 0
VFORCE__Cin_1 CIN GND DC 1.8
VFORCE__IN2 IN2 GND DC 1.8

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT TRAN V(S) V(S1)

* --- Params
.TEMP 27.0

* ELDO netlist generated with ICnet by 'vlsi' on Sat Oct 28 2017 at 04:09:33

.CONNECT GND 0

*
* Globals.
*
.global VDD GND


*
* Component pathname : $ADK/technology/ic/symbols/rxfer [SPICE]
*
*       .include /home/simulator/mentor/Library/ADK/technology/ic/symbols/rxfer/asim_lib/rxfer


*
* Component pathname : $ADK/technology/ic/symbols/prxfer [SPICE]
*
*       .include /home/simulator/mentor/Library/ADK/technology/ic/symbols/prxfer/asim_lib/prxfer

*
* Component pathname : $ADK/technology/ic/symbols/pmos4
*
.subckt PMOS4  B D G S

        X_I$410 D G S prxfer
.ends PMOS4

*
* Component pathname : $ADK/technology/ic/symbols/nmos4
*
.subckt NMOS4  B S D G

        X_I$409 D G S rxfer
.ends NMOS4

*
* MAIN CELL: Component pathname : /home/vlsi/g4/dhall_flip
*
        X_MP3 VDD N$10 N_CLK_ESC1 N$7 PMOS4
        X_MN3 GND N$7 N$10 CLK NMOS4
        X_MP2 VDD N$2 CLK N$7 PMOS4
        X_MN2 GND N$7 N$2 N_CLK_ESC1 NMOS4
        X_MP1 VDD N$2 D VDD PMOS4
        X_MN1 GND GND N$2 D NMOS4
        X_MP10 VDD OUT N$21 VDD PMOS4
        X_MN10 GND GND OUT N$21 NMOS4
        X_MP9 VDD N$24 OUT VDD PMOS4
        X_MN9 GND GND N$24 OUT NMOS4
        X_MP4 VDD N$10 N$12 VDD PMOS4
        X_MN4 GND GND N$10 N$12 NMOS4
        X_MP8 VDD N$24 CLK N$21 PMOS4
        X_MN8 GND N$21 N$24 N_CLK_ESC1 NMOS4
        X_MP7 VDD N$17 N_CLK_ESC1 N$21 PMOS4
        X_MN7 GND N$21 N$17 CLK NMOS4
        X_MP6 VDD N$17 N$12 VDD PMOS4
        X_MN6 GND GND N$17 N$12 NMOS4
        X_MP5 VDD N$12 N$7 VDD PMOS4
        X_MN5 GND GND N$12 N$7 NMOS4
*
.end

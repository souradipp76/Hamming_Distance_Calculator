* ELDO netlist generated with ICnet by 'vlsi' on Tue Oct  3 2017 at 03:27:11

.CONNECT GND 0

*
* Component pathname : /home/vlsi/dff/inverter.cir
*
.subckt INVERTER_CIR_ESC1  OUT GND IN VDD

        MN1 OUT IN GND VSS n L=1.8e-07 W=1.9e-07
        MP1 OUT IN VDD VDD p L=1.8e-07 W=1.31e-06
.ends INVERTER_CIR_ESC1

*
* MAIN CELL: Component pathname : /home/vlsi/dff/dflipflop.cir
*
        X_INVERTER_CIR4_ESC2 N$40 GND CLK VDD INVERTER_CIR_ESC1
        MN2 N$11 CLK N$24 VSS n L=1.8e-07 W=1.9e-07
        MP2 N$11 N$40 N$24 VDD p L=1.8e-07 W=1.31e-06
        MN1 N$3 N$40 N$24 VSS n L=1.8e-07 W=1.9e-07
        MP1 N$3 CLK N$24 VDD p L=1.8e-07 W=1.31e-06
        X_INVERTER_CIR3_ESC3 N$11 GND D VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR2_ESC4 OUT GND N$24 VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR1_ESC5 N$3 GND OUT VDD INVERTER_CIR_ESC1
*
.end

* Component: /home/vlsi/g4/multi Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/multi/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0.0 2000n 0

* --- Forces
VFORCE__IN IN GND DC 1.8
VFORCE__GND GND GND DC 0
VFORCE__VDD VDD GND DC 1.8
VFORCE__SEL SEL GND DC 0
VFORCE__CLK CLK GND PULSE (0 1.8 4n 1n 1n 45n 100n)
VFORCE__NCLK NCLK GND PULSE (1.8 0 4n 1n 1n 45n 100n)

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT TRAN V(O5) V(O3) V(O4) V(O2) V(O1) V(O0)

* --- Params
.TEMP 27.0

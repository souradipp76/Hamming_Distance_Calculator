* SPICE NETLIST
***************************************

.SUBCKT exclay IN2 IN1 OUT VDD GND
** N=6 EP=5 IP=0 FDC=6
M0 OUT IN2 2 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-23950 $Y=-12300 $D=1
M1 IN2 2 OUT GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-600 $Y=-12200 $D=1
M2 GND IN1 2 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=22400 $Y=-12300 $D=1
M3 OUT IN2 IN1 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-23950 $Y=5050 $D=0
M4 IN2 IN1 OUT VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-600 $Y=5150 $D=0
M5 VDD IN1 2 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=22400 $Y=5050 $D=0
.ENDS
***************************************

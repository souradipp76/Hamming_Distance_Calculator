* SPICE NETLIST
***************************************

.SUBCKT dhalllay D Clk ~Clk Out Gnd Vdd
** N=13 EP=6 IP=0 FDC=20
M0 7 D Gnd Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=157550 $Y=-5850 $D=1
M1 5 ~Clk 7 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=179650 $Y=-5850 $D=1
M2 5 Clk 8 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=204200 $Y=-5950 $D=1
M3 9 5 Gnd Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=226250 $Y=-6000 $D=1
M4 8 9 Gnd Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=248500 $Y=-6000 $D=1
M5 10 9 Gnd Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=270750 $Y=-6000 $D=1
M6 6 Clk 10 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=292850 $Y=-6000 $D=1
M7 6 ~Clk 11 Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=317400 $Y=-6100 $D=1
M8 Out 6 Gnd Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=339450 $Y=-6150 $D=1
M9 11 Out Gnd Gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=361700 $Y=-6150 $D=1
M10 7 D Vdd Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=157550 $Y=15550 $D=0
M11 5 ~Clk 8 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=179650 $Y=15550 $D=0
M12 5 Clk 7 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=204200 $Y=15450 $D=0
M13 9 5 Vdd Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=226250 $Y=15400 $D=0
M14 8 9 Vdd Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=248500 $Y=15400 $D=0
M15 10 9 Vdd Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=270750 $Y=15400 $D=0
M16 6 Clk 11 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=292850 $Y=15400 $D=0
M17 6 ~Clk 10 Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=317400 $Y=15300 $D=0
M18 Out 6 Vdd Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=339450 $Y=15250 $D=0
M19 11 Out Vdd Vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=361700 $Y=15250 $D=0
.ENDS
***************************************

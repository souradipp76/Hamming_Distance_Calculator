* ELDO netlist generated with ICnet by 'vlsi' on Thu Oct 19 2017 at 01:09:12

.CONNECT GND 0

*
* MAIN CELL: Component pathname : /home/vlsi/g4/or
*
        MN3 OUT N$7 GND VSS n L=1.8e-07 W=3.6e-07
        MP3 OUT N$7 VDD VDD p L=1.8e-07 W=1.26e-06
        MN2 N$7 IN2 GND VSS n L=1.8e-07 W=3.6e-07
        MN1 N$7 IN1 GND VSS n L=1.8e-07 W=3.6e-07
        MP2 N$5 IN1 VDD VDD p L=1.8e-07 W=2.52e-06
        MP1 N$7 IN2 N$5 VDD p L=1.8e-07 W=2.52e-06
*
.end

* File: hamminglay_pex.sp
* Created: Sat Nov  4 18:09:15 2017
* Program "Calibre xRC"
* Version "v2013.4_37.29"
* 
.include "hamminglay_pex.sp.pex"
.subckt HAMMINGLAY  CLK S1 IN1 IN2 S0
* 
* S0	S0
* IN2	IN2
* IN1	IN1
* S1	S1
* CLK	CLK
M0 N_6_M0_d N_14_M0_g N_8_M0_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M1 N_8_M1_d N_6_M1_g N_14_M1_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M2 N_23_M2_d N_6_M2_g N_14_M2_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M3 N_11_M3_d N_6_M3_g N_13_M3_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M4 N_23_M4_d N_6_M4_g N_13_M4_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M5 N_22_M5_d N_11_M5_g N_23_M5_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M6 N_23_M6_d N_22_M6_g N_12_M6_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M7 N_12_M7_d N_9_M7_g N_23_M7_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07 AD=2.349e-13
+ AS=2.349e-13
M8 N_S1_M8_d N_12_M8_g N_23_M8_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M9 N_23_M9_d N_CLK_M9_g N_7_M9_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M10 N_17_M10_d N_IN2_M10_g N_23_M10_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M11 N_17_M11_d N_IN1_M11_g N_15_M11_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M12 N_15_M12_d N_17_M12_g N_IN1_M12_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M13 N_9_M13_d N_19_M13_g N_23_M13_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M14 N_23_M14_d N_8_M14_g N_16_M14_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M15 N_19_M15_d N_10_M15_g N_16_M15_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M16 N_S0_M16_d N_8_M16_g N_18_M16_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M17 N_23_M17_d N_10_M17_g N_18_M17_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M18 N_8_M18_d N_18_M18_g N_S0_M18_s N_23_X40.M0_b n L=1.8e-07 W=3.6e-07
+ AD=2.349e-13 AS=2.349e-13
M19 N_6_M19_d N_6_M19_g N_8_M19_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M20 N_8_M20_d N_6_M20_g N_6_M20_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M21 N_21_M21_d N_6_M21_g N_14_M21_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M22 N_11_M22_d N_6_M22_g N_21_M22_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M23 N_21_M23_d N_6_M23_g N_11_M23_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M24 N_22_M24_d N_11_M24_g N_21_M24_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M25 N_20_M25_d N_22_M25_g N_21_M25_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M26 N_12_M26_d N_9_M26_g N_20_M26_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M27 N_S1_M27_d N_12_M27_g N_21_M27_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M28 N_21_M28_d N_CLK_M28_g N_7_M28_s N_21_X40.M30_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M29 N_17_M29_d N_IN2_M29_g N_24_M29_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M30 N_IN2_M30_d N_IN1_M30_g N_15_M30_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M31 N_15_M31_d N_IN2_M31_g N_IN1_M31_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M32 N_9_M32_d N_19_M32_g N_24_M32_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M33 N_24_M33_d N_8_M33_g N_19_M33_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M34 N_19_M34_d N_10_M34_g N_24_M34_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M35 N_S0_M35_d N_8_M35_g N_10_M35_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M36 N_24_M36_d N_10_M36_g N_18_M36_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
M37 N_8_M37_d N_10_M37_g N_S0_M37_s N_24_M29_b p L=1.8e-07 W=1.26e-06
+ AD=6.237e-13 AS=6.237e-13
mX40.M0 N_X40.14_X40.M0_d N_15_X40.M0_g N_23_X40.M0_s N_23_X40.M0_b n L=1.8e-07
+ W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M1 N_X40.15_X40.M1_d N_6_X40.M1_g N_23_X40.M1_s N_23_X40.M0_b n L=1.8e-07
+ W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M2 N_X40.16_X40.M2_d N_6_X40.M2_g N_23_X40.M2_s N_23_X40.M0_b n L=1.8e-07
+ W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M3 N_X40.8_X40.M3_d N_7_X40.M3_g N_X40.14_X40.M3_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M4 N_X40.9_X40.M4_d N_7_X40.M4_g N_X40.15_X40.M4_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M5 N_X40.10_X40.M5_d N_7_X40.M5_g N_X40.16_X40.M5_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M6 N_X40.8_X40.M6_d N_CLK_X40.M6_g N_X40.17_X40.M6_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M7 N_X40.9_X40.M7_d N_CLK_X40.M7_g N_X40.18_X40.M7_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M8 N_X40.10_X40.M8_d N_CLK_X40.M8_g N_X40.19_X40.M8_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M9 N_X40.20_X40.M9_d N_X40.8_X40.M9_g N_23_X40.M9_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M10 N_X40.21_X40.M10_d N_X40.9_X40.M10_g N_23_X40.M10_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M11 N_X40.22_X40.M11_d N_X40.10_X40.M11_g N_23_X40.M11_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M12 N_X40.17_X40.M12_d N_X40.20_X40.M12_g N_23_X40.M12_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M13 N_X40.18_X40.M13_d N_X40.21_X40.M13_g N_23_X40.M13_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M14 N_X40.19_X40.M14_d N_X40.22_X40.M14_g N_23_X40.M14_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M15 N_X40.23_X40.M15_d N_X40.20_X40.M15_g N_23_X40.M15_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M16 N_X40.24_X40.M16_d N_X40.21_X40.M16_g N_23_X40.M16_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M17 N_X40.25_X40.M17_d N_X40.22_X40.M17_g N_23_X40.M17_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M18 N_X40.11_X40.M18_d N_CLK_X40.M18_g N_X40.23_X40.M18_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M19 N_X40.12_X40.M19_d N_CLK_X40.M19_g N_X40.24_X40.M19_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M20 N_X40.13_X40.M20_d N_CLK_X40.M20_g N_X40.25_X40.M20_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M21 N_X40.11_X40.M21_d N_7_X40.M21_g N_X40.26_X40.M21_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M22 N_X40.12_X40.M22_d N_7_X40.M22_g N_X40.27_X40.M22_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M23 N_X40.13_X40.M23_d N_7_X40.M23_g N_X40.28_X40.M23_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M24 N_6_X40.M24_d N_X40.11_X40.M24_g N_23_X40.M24_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M25 N_6_X40.M25_d N_X40.12_X40.M25_g N_23_X40.M25_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M26 N_10_X40.M26_d N_X40.13_X40.M26_g N_23_X40.M26_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M27 N_X40.26_X40.M27_d N_6_X40.M27_g N_23_X40.M27_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M28 N_X40.27_X40.M28_d N_6_X40.M28_g N_23_X40.M28_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M29 N_X40.28_X40.M29_d N_10_X40.M29_g N_23_X40.M29_s N_23_X40.M0_b n
+ L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13
mX40.M30 N_X40.14_X40.M30_d N_15_X40.M30_g N_21_X40.M30_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M31 N_X40.15_X40.M31_d N_6_X40.M31_g N_21_X40.M31_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M32 N_X40.16_X40.M32_d N_6_X40.M32_g N_21_X40.M32_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M33 N_X40.8_X40.M33_d N_7_X40.M33_g N_X40.17_X40.M33_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M34 N_X40.9_X40.M34_d N_7_X40.M34_g N_X40.18_X40.M34_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M35 N_X40.10_X40.M35_d N_7_X40.M35_g N_X40.19_X40.M35_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M36 N_X40.8_X40.M36_d N_CLK_X40.M36_g N_X40.14_X40.M36_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M37 N_X40.9_X40.M37_d N_CLK_X40.M37_g N_X40.15_X40.M37_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M38 N_X40.10_X40.M38_d N_CLK_X40.M38_g N_X40.16_X40.M38_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M39 N_X40.20_X40.M39_d N_X40.8_X40.M39_g N_21_X40.M39_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M40 N_X40.21_X40.M40_d N_X40.9_X40.M40_g N_21_X40.M40_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M41 N_X40.22_X40.M41_d N_X40.10_X40.M41_g N_21_X40.M41_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M42 N_X40.17_X40.M42_d N_X40.20_X40.M42_g N_21_X40.M42_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M43 N_X40.18_X40.M43_d N_X40.21_X40.M43_g N_21_X40.M43_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M44 N_X40.19_X40.M44_d N_X40.22_X40.M44_g N_21_X40.M44_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M45 N_X40.23_X40.M45_d N_X40.20_X40.M45_g N_21_X40.M45_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M46 N_X40.24_X40.M46_d N_X40.21_X40.M46_g N_21_X40.M46_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M47 N_X40.25_X40.M47_d N_X40.22_X40.M47_g N_21_X40.M47_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M48 N_X40.11_X40.M48_d N_CLK_X40.M48_g N_X40.26_X40.M48_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M49 N_X40.12_X40.M49_d N_CLK_X40.M49_g N_X40.27_X40.M49_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M50 N_X40.13_X40.M50_d N_CLK_X40.M50_g N_X40.28_X40.M50_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M51 N_X40.11_X40.M51_d N_7_X40.M51_g N_X40.23_X40.M51_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M52 N_X40.12_X40.M52_d N_7_X40.M52_g N_X40.24_X40.M52_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M53 N_X40.13_X40.M53_d N_7_X40.M53_g N_X40.25_X40.M53_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M54 N_6_X40.M54_d N_X40.11_X40.M54_g N_21_X40.M54_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M55 N_6_X40.M55_d N_X40.12_X40.M55_g N_21_X40.M55_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M56 N_10_X40.M56_d N_X40.13_X40.M56_g N_21_X40.M56_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M57 N_X40.26_X40.M57_d N_6_X40.M57_g N_21_X40.M57_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M58 N_X40.27_X40.M58_d N_6_X40.M58_g N_21_X40.M58_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
mX40.M59 N_X40.28_X40.M59_d N_10_X40.M59_g N_21_X40.M59_s N_21_X40.M30_b p
+ L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13
*
.include "hamminglay_pex.sp.HAMMINGLAY.pxi"
*
.ends
*
*

* Component: /home/vlsi/dff/inverter.cir Viewpoint: tsmc018a

.INCLUDE /home/vlsi/dff/inverter.cir/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0.0 100n 0 UIC

* --- Forces
VFORCE___VDD VDD GND DC 1.8
VFORCE___GND GND GND DC 0
VFORCE__IN IN GND PULSE (0 1.8 0n 1n 1n 25n 50n)

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PROBE TRAN V(OUT)

* --- Params
.TEMP 27.0

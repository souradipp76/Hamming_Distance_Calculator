* SPICE NETLIST
***************************************

.SUBCKT nwell_contact
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT halfaddlay IN1 IN2 S GND VDD C
** N=9 EP=6 IP=2 FDC=12
M0 S IN2 3 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-23950 $Y=-12300 $D=1
M1 IN2 3 S GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=-600 $Y=-12200 $D=1
M2 GND IN1 3 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=22400 $Y=-12300 $D=1
M3 5 IN1 4 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=44550 $Y=-12350 $D=1
M4 GND IN2 4 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=66600 $Y=-12450 $D=1
M5 C 5 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=88900 $Y=-12500 $D=1
M6 S IN2 IN1 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-23950 $Y=5050 $D=0
M7 IN2 IN1 S VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=-600 $Y=5150 $D=0
M8 VDD IN1 3 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=22400 $Y=5050 $D=0
M9 5 IN1 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=44550 $Y=5000 $D=0
M10 VDD IN2 5 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=66600 $Y=4900 $D=0
M11 C 5 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=88900 $Y=4850 $D=0
.ENDS
***************************************

* ELDO netlist generated with ICnet by 'vlsi' on Mon Oct  9 2017 at 00:22:06

.CONNECT GND 0

*
* MAIN CELL: Component pathname : /home/vlsi/dff/inverter.cir
*
.SUBCKT invstage1_lay OUT IN GND VDD 
        MN1 OUT IN GND GND n L=1.8e-07 W=1.9e-07
        MP1 OUT IN VDD VDD p L=1.8e-07 W=1.31e-06
*
.ends




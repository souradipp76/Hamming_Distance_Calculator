* Component: /home/vlsi/dff/sipopiso.cir Viewpoint: tsmc018a

.INCLUDE /home/vlsi/dff/sipopiso.cir/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000.0
.OPTION NOASCII

* - Analysis Setup - DCOP
.OPTION PROBEOP2
.OP

* - Analysis Setup - Trans
.TRAN 0.0 100n 0 UIC

* --- Forces
VFORCE__A A GND DC 0
VFORCE__B B GND DC 0
VFORCE__C C GND DC 0
VFORCE__D D GND DC 0
VFORCE__GND GND GND DC 0
VFORCE__S S GND DC 0
VFORCE__VDD VDD GND DC 1.8
VFORCE__SIN SIN GND PATTERN 1.8 0 0 1n 1n 50n 1101 R=-1
VFORCE__CLK CLK GND PATTERN 1.8 0 25n 1n 1n 50n 1010 R=-1

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT DC V(SO)
.PLOT TRAN V(SO)

* --- Params
.TEMP 27.0

* SPICE NETLIST
***************************************

.SUBCKT nwell_contact
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sipo2 1 2 3 4 5 gnd vdd
** N=28 EP=7 IP=2 FDC=60
* PORT gnd gnd 261000 -24225 METAL1
* PORT vdd vdd 261400 50825 METAL1
* PORT gnd gnd 258900 -169225 METAL1
* PORT vdd vdd 259000 -95375 METAL1
M0 14 5 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=157550 $Y=-5850 $D=1
M1 15 4 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=157850 $Y=-42900 $D=1
M2 16 4 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=158050 $Y=-152250 $D=1
M3 8 2 14 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=179650 $Y=-5850 $D=1
M4 9 2 15 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=179950 $Y=-42900 $D=1
M5 10 2 16 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=180150 $Y=-152250 $D=1
M6 8 1 17 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=204200 $Y=-5950 $D=1
M7 9 1 18 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=204500 $Y=-42800 $D=1
M8 10 1 19 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=204700 $Y=-152350 $D=1
M9 20 8 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=226250 $Y=-6000 $D=1
M10 21 9 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=226550 $Y=-42750 $D=1
M11 22 10 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=226750 $Y=-152400 $D=1
M12 17 20 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=248500 $Y=-6000 $D=1
M13 18 21 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=248800 $Y=-42750 $D=1
M14 19 22 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=249000 $Y=-152400 $D=1
M15 23 20 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=270750 $Y=-6000 $D=1
M16 24 21 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=271050 $Y=-42750 $D=1
M17 25 22 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=271250 $Y=-152400 $D=1
M18 11 1 23 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=292850 $Y=-6000 $D=1
M19 12 1 24 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=293150 $Y=-42750 $D=1
M20 13 1 25 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=293350 $Y=-152400 $D=1
M21 11 2 26 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=317400 $Y=-6100 $D=1
M22 12 2 27 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=317700 $Y=-42650 $D=1
M23 13 2 28 gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=317900 $Y=-152500 $D=1
M24 4 11 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=339450 $Y=-6150 $D=1
M25 4 12 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=339750 $Y=-42600 $D=1
M26 3 13 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=339950 $Y=-152550 $D=1
M27 26 4 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=361700 $Y=-6150 $D=1
M28 27 4 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=362000 $Y=-42600 $D=1
M29 28 3 gnd gnd N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=362200 $Y=-152550 $D=1
M30 14 5 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=157550 $Y=15550 $D=0
M31 15 4 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=157850 $Y=-74300 $D=0
M32 16 4 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=158050 $Y=-130850 $D=0
M33 8 2 17 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=179650 $Y=15550 $D=0
M34 9 2 18 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=179950 $Y=-74300 $D=0
M35 10 2 19 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=180150 $Y=-130850 $D=0
M36 8 1 14 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=204200 $Y=15450 $D=0
M37 9 1 15 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=204500 $Y=-74200 $D=0
M38 10 1 16 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=204700 $Y=-130950 $D=0
M39 20 8 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=226250 $Y=15400 $D=0
M40 21 9 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=226550 $Y=-74150 $D=0
M41 22 10 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=226750 $Y=-131000 $D=0
M42 17 20 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=248500 $Y=15400 $D=0
M43 18 21 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=248800 $Y=-74150 $D=0
M44 19 22 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=249000 $Y=-131000 $D=0
M45 23 20 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=270750 $Y=15400 $D=0
M46 24 21 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=271050 $Y=-74150 $D=0
M47 25 22 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=271250 $Y=-131000 $D=0
M48 11 1 26 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=292850 $Y=15400 $D=0
M49 12 1 27 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=293150 $Y=-74150 $D=0
M50 13 1 28 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=293350 $Y=-131000 $D=0
M51 11 2 23 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=317400 $Y=15300 $D=0
M52 12 2 24 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=317700 $Y=-74050 $D=0
M53 13 2 25 vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=317900 $Y=-131100 $D=0
M54 4 11 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=339450 $Y=15250 $D=0
M55 4 12 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=339750 $Y=-74000 $D=0
M56 3 13 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=339950 $Y=-131150 $D=0
M57 26 4 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=361700 $Y=15250 $D=0
M58 27 4 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=362000 $Y=-74000 $D=0
M59 28 3 vdd vdd P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=362200 $Y=-131150 $D=0
.ENDS
***************************************
.SUBCKT hamminglay clk s1 in1 in2 s0
** N=24 EP=5 IP=9 FDC=98
* PORT clk clk 444350 345050 METAL4
* PORT s1 s1 538950 312950 METAL4
* PORT in1 in1 494900 342400 METAL4
* PORT in2 in2 518400 342750 METAL4
* PORT s0 s0 535350 131300 METAL4
M0 6 14 8 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451150 $Y=136500 $D=1
M1 8 6 14 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451250 $Y=113150 $D=1
M2 23 6 14 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451250 $Y=159500 $D=1
M3 11 6 13 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451300 $Y=181650 $D=1
M4 23 6 13 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451400 $Y=203700 $D=1
M5 22 11 23 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451450 $Y=226000 $D=1
M6 23 22 12 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451500 $Y=248200 $D=1
M7 12 9 23 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451550 $Y=271600 $D=1
M8 s1 12 23 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451550 $Y=294500 $D=1
M9 23 clk 7 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451750 $Y=328400 $D=1
M10 17 in2 23 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=482800 $Y=248850 $D=1
M11 17 in1 15 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=482800 $Y=295200 $D=1
M12 15 17 in1 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=482900 $Y=271850 $D=1
M13 9 19 23 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483000 $Y=225750 $D=1
M14 23 8 16 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483050 $Y=203450 $D=1
M15 19 10 16 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483150 $Y=181400 $D=1
M16 s0 8 18 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483200 $Y=112900 $D=1
M17 23 10 18 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483200 $Y=159250 $D=1
M18 8 18 s0 23 N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483300 $Y=136250 $D=1
M19 6 6 8 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=423800 $Y=136500 $D=0
M20 8 6 6 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=423900 $Y=113150 $D=0
M21 21 6 14 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=423900 $Y=159500 $D=0
M22 11 6 21 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=423950 $Y=181650 $D=0
M23 21 6 11 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424050 $Y=203700 $D=0
M24 22 11 21 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424100 $Y=226000 $D=0
M25 20 22 21 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424150 $Y=248200 $D=0
M26 12 9 20 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424200 $Y=271600 $D=0
M27 s1 12 21 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424200 $Y=294500 $D=0
M28 21 clk 7 21 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424250 $Y=328400 $D=0
M29 17 in2 24 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500150 $Y=248850 $D=0
M30 in2 in1 15 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500150 $Y=295200 $D=0
M31 15 in2 in1 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500250 $Y=271850 $D=0
M32 9 19 24 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500350 $Y=225750 $D=0
M33 24 8 19 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500400 $Y=203450 $D=0
M34 19 10 24 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500500 $Y=181400 $D=0
M35 s0 8 10 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500550 $Y=112900 $D=0
M36 24 10 18 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500550 $Y=159250 $D=0
M37 8 10 s0 24 P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500650 $Y=136250 $D=0
X40 clk 7 10 6 15 23 21 sipo2 $T=540300 279250 1 180 $X=160850 $Y=104250
.ENDS
***************************************

* Component: /home/vlsi/g4/inv Viewpoint: tsmc018a

.INCLUDE /home/vlsi/g4/inv/tsmc018a/netlist.spi
.INCLUDE $ADK/technology/ic/models/tsmc018.mod
.OPTION AEX
.OPTION ENGNOT
.OPTION LIMPROBE=10000
.OPTION NOASCII

* - Analysis Setup - Trans
.TRAN 0 100n 0

* --- Forces
VFORCE__IN IN GND PULSE (0 1.8 0 1n 1n 20n 50n)
VFORCE__GND GND GND DC 0
VFORCE__VDD VDD GND DC 1.8

* --- Global Outputs
.PROBE V SG

* --- Waveform Outputs
.PLOT TRAN V(IN) V(OUT)

* --- Params
.TEMP 27

* ELDO netlist generated with ICnet by 'vlsi' on Sat Oct 28 2017 at 02:03:46

.CONNECT GND 0

*
* Component pathname : /home/vlsi/dff/inverter.cir
*
.subckt INVERTER_CIR_ESC1  OUT GND IN VDD

        MN1 OUT IN GND VSS n L=1.8e-07 W=1.9e-07
        MP1 OUT IN VDD VDD p L=1.8e-07 W=1.31e-06
.ends INVERTER_CIR_ESC1

*
* Component pathname : /home/vlsi/dff/Dflipflopnoinvnew.cir
*
.subckt DFLIPFLOPNOINVNEW_CIR_ESC2  OUT CLK D GND NCLK VDD

        MN2 N$7 CLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP2 N$7 NCLK N$56 VDD p L=1.8e-07 W=1.31e-06
        MN1 N$4 NCLK N$56 VSS n L=1.8e-07 W=1.9e-07
        MP1 N$4 CLK N$56 VDD p L=1.8e-07 W=1.31e-06
        X_INVERTER_CIR3_ESC3 OUT GND N$56 VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR2_ESC4 N$7 GND D VDD INVERTER_CIR_ESC1
        X_INVERTER_CIR1_ESC5 N$4 GND OUT VDD INVERTER_CIR_ESC1
.ends DFLIPFLOPNOINVNEW_CIR_ESC2

*
* Component pathname : /home/vlsi/dff/masterslaveDflipflopnew.cir
*
.subckt MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6  OUT CLEAR CLK D GND NCLK PRESET
+ VDD

        X_DFLIPFLOPNOINVNEW_CIR1_ESC7 N$34 NCLK D GND CLK VDD DFLIPFLOPNOINVNEW_CIR_ESC2
        X_DFLIPFLOPNOINVNEW_CIR2_ESC8 OUT CLK N$34 GND NCLK VDD DFLIPFLOPNOINVNEW_CIR_ESC2
.ends MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6

*
* MAIN CELL: Component pathname : /home/vlsi/g4/sipo.cir
*
        X_DFF3 P3 N$45 CLK P2 GND NCLK N$44 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_DFF2 P2 N$45 CLK P1 GND NCLK N$44 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
        X_DFF1 P1 N$45 CLK SIN GND NCLK N$44 VDD MASTERSLAVEDFLIPFLOPNEW_CIR_ESC6
*
.end

* ELDO netlist generated with ICnet by 'vlsi' on Mon Oct  9 2017 at 08:12:44

.CONNECT GND 0

*
* MAIN CELL: Component pathname : /home/vlsi/dff/inverter.cir
*
        MN1 OUT IN GND VSS n L=1.8e-07 W=1.9e-07
        MP1 OUT IN VDD VDD p L=1.8e-07 W=1.31e-06
*
.end

* ELDO netlist generated with ICnet by 'vlsi' on Tue Oct 24 2017 at 10:05:05

.CONNECT GND 0

*
* MAIN CELL: Component pathname : /home/vlsi/g4/xor
*
        MN7 OUT N$22 GND VSS n L=1.8e-07 W=3.6e-07
        MP7 OUT N$22 VDD VDD p L=1.8e-07 W=1.26e-06
        MP6 IN2N IN2 VDD VDD p L=1.8e-07 W=1.26e-06
        MN6 IN2N IN2 GND VSS n L=1.8e-07 W=3.6e-07
        MP5 INN IN1 VDD VDD p L=1.8e-07 W=1.26e-06
        MN5 INN IN1 GND VSS n L=1.8e-07 W=3.6e-07
        MN1 N$22 INN N$24 VSS n L=1.8e-07 W=7.2e-07
        MN4 N$2 IN2N GND VSS n L=1.8e-07 W=7.2e-07
        MN3 N$24 IN2 GND VSS n L=1.8e-07 W=7.2e-07
        MN2 N$22 IN1 N$2 VSS n L=1.8e-07 W=7.2e-07
        MP4 N$22 IN2N N$7 VDD p L=1.8e-07 W=2.52e-06
        MP3 N$7 INN VDD VDD p L=1.8e-07 W=2.52e-06
        MP2 N$22 IN2 N$31 VDD p L=1.8e-07 W=2.52e-06
        MP1 N$31 IN1 VDD VDD p L=1.8e-07 W=2.52e-06
*
.end

* SPICE NETLIST
***************************************

.SUBCKT nwell_contact
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT hamming_lay clk s1 in2 in1 s0 VDD GND
** N=45 EP=7 IP=4 FDC=98
M0 GND 1 18 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=176050 $Y=126750 $D=1
M1 GND 3 19 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=176250 $Y=236700 $D=1
M2 GND 15 20 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=176550 $Y=273150 $D=1
M3 GND 9 1 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=198300 $Y=126750 $D=1
M4 GND 10 3 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=198500 $Y=236700 $D=1
M5 GND 11 15 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=198800 $Y=273150 $D=1
M6 18 2 9 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=220350 $Y=126800 $D=1
M7 19 2 10 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=220550 $Y=236650 $D=1
M8 20 2 11 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=220850 $Y=273200 $D=1
M9 21 clk 9 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=244900 $Y=126900 $D=1
M10 22 clk 10 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=245100 $Y=236550 $D=1
M11 23 clk 11 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=245400 $Y=273300 $D=1
M12 GND 24 21 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=267000 $Y=126900 $D=1
M13 GND 25 22 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=267200 $Y=236550 $D=1
M14 GND 26 23 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=267500 $Y=273300 $D=1
M15 GND 24 27 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=289250 $Y=126900 $D=1
M16 GND 25 28 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=289450 $Y=236550 $D=1
M17 GND 26 29 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=289750 $Y=273300 $D=1
M18 GND 12 24 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=311500 $Y=126900 $D=1
M19 GND 13 25 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=311700 $Y=236550 $D=1
M20 GND 14 26 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=312000 $Y=273300 $D=1
M21 27 clk 12 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=333550 $Y=126950 $D=1
M22 28 clk 13 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=333750 $Y=236500 $D=1
M23 29 clk 14 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=334050 $Y=273350 $D=1
M24 30 2 12 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=358100 $Y=127050 $D=1
M25 31 2 13 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=358300 $Y=236400 $D=1
M26 32 2 14 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=358600 $Y=273450 $D=1
M27 GND 3 30 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=380200 $Y=127050 $D=1
M28 GND 15 31 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=380400 $Y=236400 $D=1
M29 GND 37 32 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=380700 $Y=273450 $D=1
M30 3 36 16 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451150 $Y=136500 $D=1
M31 16 3 36 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451250 $Y=113150 $D=1
M32 GND 15 36 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451250 $Y=159500 $D=1
M33 33 15 35 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451300 $Y=181650 $D=1
M34 GND 3 35 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451400 $Y=203700 $D=1
M35 45 33 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451450 $Y=226000 $D=1
M36 GND 45 34 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451500 $Y=248200 $D=1
M37 34 17 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451550 $Y=271600 $D=1
M38 s1 34 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451550 $Y=294500 $D=1
M39 GND clk 2 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=451650 $Y=328700 $D=1
M40 39 in1 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=482800 $Y=248850 $D=1
M41 39 in2 37 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=482800 $Y=295200 $D=1
M42 37 39 in2 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=482900 $Y=271850 $D=1
M43 17 41 GND GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483000 $Y=225750 $D=1
M44 GND 16 38 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483050 $Y=203450 $D=1
M45 41 1 38 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483150 $Y=181400 $D=1
M46 s0 16 40 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483200 $Y=112900 $D=1
M47 GND 1 40 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483200 $Y=159250 $D=1
M48 16 40 s0 GND N L=1.8e-07 W=3.6e-07 AD=2.349e-13 AS=2.349e-13 $X=483300 $Y=136250 $D=1
M49 VDD 1 18 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=176050 $Y=148150 $D=0
M50 VDD 3 19 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=176250 $Y=205300 $D=0
M51 VDD 15 20 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=176550 $Y=294550 $D=0
M52 VDD 9 1 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=198300 $Y=148150 $D=0
M53 VDD 10 3 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=198500 $Y=205300 $D=0
M54 VDD 11 15 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=198800 $Y=294550 $D=0
M55 21 2 9 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=220350 $Y=148200 $D=0
M56 22 2 10 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=220550 $Y=205250 $D=0
M57 23 2 11 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=220850 $Y=294600 $D=0
M58 18 clk 9 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=244900 $Y=148300 $D=0
M59 19 clk 10 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=245100 $Y=205150 $D=0
M60 20 clk 11 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=245400 $Y=294700 $D=0
M61 VDD 24 21 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=267000 $Y=148300 $D=0
M62 VDD 25 22 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=267200 $Y=205150 $D=0
M63 VDD 26 23 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=267500 $Y=294700 $D=0
M64 VDD 24 27 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=289250 $Y=148300 $D=0
M65 VDD 25 28 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=289450 $Y=205150 $D=0
M66 VDD 26 29 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=289750 $Y=294700 $D=0
M67 VDD 12 24 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=311500 $Y=148300 $D=0
M68 VDD 13 25 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=311700 $Y=205150 $D=0
M69 VDD 14 26 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=312000 $Y=294700 $D=0
M70 30 clk 12 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=333550 $Y=148350 $D=0
M71 31 clk 13 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=333750 $Y=205100 $D=0
M72 32 clk 14 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=334050 $Y=294750 $D=0
M73 27 2 12 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=358100 $Y=148450 $D=0
M74 28 2 13 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=358300 $Y=205000 $D=0
M75 29 2 14 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=358600 $Y=294850 $D=0
M76 VDD 3 30 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=380200 $Y=148450 $D=0
M77 VDD 15 31 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=380400 $Y=205000 $D=0
M78 VDD 37 32 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=380700 $Y=294850 $D=0
M79 3 15 16 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=423800 $Y=136500 $D=0
M80 16 3 15 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=423900 $Y=113150 $D=0
M81 VDD 15 36 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=423900 $Y=159500 $D=0
M82 33 15 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=423950 $Y=181650 $D=0
M83 VDD 3 33 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424050 $Y=203700 $D=0
M84 45 33 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424100 $Y=226000 $D=0
M85 44 45 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424150 $Y=248200 $D=0
M86 VDD clk 2 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424150 $Y=328700 $D=0
M87 34 17 44 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424200 $Y=271600 $D=0
M88 s1 34 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=424200 $Y=294500 $D=0
M89 39 in1 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500150 $Y=248850 $D=0
M90 in1 in2 37 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500150 $Y=295200 $D=0
M91 37 in1 in2 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500250 $Y=271850 $D=0
M92 17 41 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500350 $Y=225750 $D=0
M93 VDD 16 41 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500400 $Y=203450 $D=0
M94 41 1 VDD VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500500 $Y=181400 $D=0
M95 s0 16 1 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500550 $Y=112900 $D=0
M96 VDD 1 40 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500550 $Y=159250 $D=0
M97 16 1 s0 VDD P L=1.8e-07 W=1.26e-06 AD=6.237e-13 AS=6.237e-13 $X=500650 $Y=136250 $D=0
.ENDS
***************************************
